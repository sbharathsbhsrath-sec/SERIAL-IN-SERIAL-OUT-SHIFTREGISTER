module siso(clk, sin, q); 
input clk; 
input sin; 
output [3:0] q; 
reg [3:0] q; 
always @(posedge clk) 
begin 
q[0] <= sin; 
q[1] <= q[0]; 
q[2] <= q[1]; 
q[3] <= q[2]; 
end 
endmodule 
